`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company:   CS141
// Engineer:  Avinash Uttamchandani
//
////////////////////////////////////////////////////////////////////////////////

`include "alu_defines.v"

module test_alu;

	// Inputs
	reg [31:0] X;
	reg [31:0] Y;
	reg [3:0] op_code;

	// Outputs
	wire [31:0] Z;
	wire equal;
	wire overflow;
	wire zero;

	// Instantiate the Unit Under Test (UUT)
	alu uut (
		.X(X), 
		.Y(Y), 
		.Z(Z), 
		.op_code(op_code), 
		.equal(equal), 
		.overflow(overflow), 
		.zero(zero)
	);

	// HINT: 'integer' variables might be useful
	
	initial begin
		op_code = `ALU_OP_AND;
		
			  X = 32'b00000000000000000000000000000000; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b11111111111111111111111111111111;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b11111111111111111111111111111111;
		
		#10; op_code = `ALU_OP_OR;
		
		     X = 32'b00000000000000000000000000000000; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b11111111111111111111111111111111;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b11111111111111111111111111111111;
		
		#10; op_code = `ALU_OP_XOR;
				
		     X = 32'b00000000000000000000000000000000; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b11111111111111111111111111111111;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b11111111111111111111111111111111;
		
		#10; op_code =`ALU_OP_NOR;
			
		     X = 32'b00000000000000000000000000000000; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b00000000000000000000000000000000; Y = 32'b11111111111111111111111111111111;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b10101010101010101010101010101010;
		#10; X = 32'b10101010101010101010101010101010; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b01010101010101010101010101010101;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b11111111111111111111111111111111;
		
		#10; op_code = `ALU_OP_ADD;
				
		     X = 32'b00000000000000000000000000000000; Y = 32'b00000000000000000000000000000000;
		#10; X = 32'b00000000000000000000000000000001; Y = 32'b00000000000000000000000000000001;
		#10; X = 32'b00000000000000000000000000000010; Y = 32'b00000000000000000000000000000001;
		#10; X = 32'b01111111111111111111111111111111; Y = 32'b00000000000000000000000000000001;
		#10; X = 32'b11111111111111111111111111111111; Y = 32'b00000000000000000000000000000001; //overflow case
		#10; X = 32'b01111111111111111111111111111111; Y = 32'b01111111111111111111111111111111;
		#10; X = 32'b01001101001011111001100111111101; Y = 32'b11100101111001000001110101101001; //1294965245 + (-438035095) = 856930150
		#10;

		
		$finish;
	
	end
	
	//a checker
	always @(X,Y,op_code) begin
		#1;
		case (op_code)
			`ALU_OP_AND : begin
				//only executes when the op code is 0000 (AND)
				if( Z !== (X & Y) ) begin
					$display("ERROR: AND:  op_code = %b, X = %h, Y = %h, Z = %h", op_code, X, Y, Z);
					//error = error + 1;
				end
			end
			// ADD IN YOUR OWN OP CODE CHECKERS HERE!!!
			`ALU_OP_XOR : begin
			end
			`ALU_OP_OR : begin
			end
			`ALU_OP_NOR: begin
			end
			`ALU_OP_ADD: begin
			end
			`ALU_OP_SUB: begin
			end
			`ALU_OP_SLT: begin
			end
			`ALU_OP_SRL: begin
			end
			`ALU_OP_SLL: begin
			end
			`ALU_OP_SRA: begin
			end
			default : begin
				//executes at default
				if (Z !== 32'd0) begin
					$display("ERROR HAPPENED! invalid op code, Z was not zero, op_code = %b, X = %h, Y = %h, Z = %h", op_code, X, Y, Z);
				end
			end
		endcase
		
	end
	
endmodule

